module token

pub const constants_tok = {
	'true': TokenType.boolean_true
	'false': TokenType.boolean_false
	'default': TokenType.boolean_default
	'on': TokenType.boolean_enable
	'off': TokenType.boolean_disable
}
