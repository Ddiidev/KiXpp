module token

pub const builtin_functions_tok = {
	'ubound': TokenType.builtin_function
}
